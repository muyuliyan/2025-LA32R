module trap_handler (
    ports
);
    
endmodule