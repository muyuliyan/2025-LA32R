module int_controler (
    ports
);
    
endmodule